`timescale 1ns/1ps
module exponential(input clock, output successful);

    (* ram_style = "distributed" *) reg [95:0] LUT [0:31];
    reg [31:0] x = 32'b11000000001100000000000000000000;
    reg [9:0] index;
    reg valid_x_l;
    reg reset;
    reg [1:0] delay;
    reg start_delaying;
    wire compared;
    wire [7:0] x_lesser_than_x_l;
    wire [31:0] e_x;
    
    floating_point_2 comparing_x_l(
      .aclk(clock),                                  // input wire aclk
      .aresetn(reset),                            // input wire aresetn
      .s_axis_a_tvalid(1),            // input wire s_axis_a_tvalid
      .s_axis_a_tready(),            // output wire s_axis_a_tready
      .s_axis_a_tdata(x),              // input wire [31 : 0] s_axis_a_tdata
      .s_axis_b_tvalid(valid_x_l),            // input wire s_axis_b_tvalid
      .s_axis_b_tready(),            // output wire s_axis_b_tready
      .s_axis_b_tdata(LUT[index][95:64]),              // input wire [31 : 0] s_axis_b_tdata
      .m_axis_result_tvalid(compared),  // output wire m_axis_result_tvalid
      .m_axis_result_tready(valid_x_l),  // input wire m_axis_result_tready
      .m_axis_result_tdata(x_lesser_than_x_l)    // output wire [7 : 0] m_axis_result_tdata
    );
    
    floating_point_1 computing_e_x(
      .aclk(clock),                                  // input wire aclk
      .s_axis_a_tvalid(x_lesser_than_x_l[0]),            // input wire s_axis_a_tvalid
      .s_axis_a_tready(),            // output wire s_axis_a_tready
      .s_axis_a_tdata(LUT[index - 10'b0000000001][63:32]),              // input wire [31 : 0] s_axis_a_tdata
      .s_axis_b_tvalid(1),            // input wire s_axis_b_tvalid
      .s_axis_b_tready(),            // output wire s_axis_b_tready
      .s_axis_b_tdata(x),              // input wire [31 : 0] s_axis_b_tdata
      .s_axis_c_tvalid(x_lesser_than_x_l[0]),            // input wire s_axis_c_tvalid
      .s_axis_c_tready(),            // output wire s_axis_c_tready
      .s_axis_c_tdata(LUT[index - 10'b0000000001][31:0]),              // input wire [31 : 0] s_axis_c_tdata
      .m_axis_result_tvalid(successful),  // output wire m_axis_result_tvalid
      .m_axis_result_tready(x_lesser_than_x_l[0]),  // input wire m_axis_result_tready
      .m_axis_result_tdata(e_x)    // output wire [31 : 0] m_axis_result_tdata
    );
    
    initial begin
        LUT[0] = 96'b110000010000000000000000000000000011100111000111110100010000001100111011010111011100110100100101;
        LUT[1] = 96'b110000001111100000000000000000000011101000000000010010001110001100111011100010100110001111110000;
        LUT[2] = 96'b110000001111000000000000000000000011101000100100101110001000100000111011101011001000110010011011;
        LUT[3] = 96'b110000001110100000000000000000000011101001010011100000010111011100111011110101101111001010110100;
        LUT[4] = 96'b110000001110000000000000000000000011101010000111110010100001010000111100000001011100000110000111;
        LUT[5] = 96'b110000001101100000000000000000000011101010101110010110110110010000111100001001100100110000100011;
        LUT[6] = 96'b110000001101000000000000000000000011101011011111111000001111101000111100010011101000100010101100;
        LUT[7] = 96'b110000001100100000000000000000000011101100001111101110111010100100111100100000000001101100010000;
        LUT[8] = 96'b110000001100000000000000000000000011101100111000100011101001000000111100100111101011100100111110;
        LUT[9] = 96'b110000001011100000000000000000000011101101101100111110011100100100111100110001000110011001001111;
        LUT[10] = 96'b110000001011000000000000000000000011101110011000001001000011010000111100111100101010110001011101;
        LUT[11] = 96'b110000001010100000000000000000000011101111000011010110100111110000111101000101011011000111001101;
        LUT[12] = 96'b110000001010000000000000000000000011101111111010110101101011110000111101001110000101111101110101;
        LUT[13] = 96'b110000001001100000000000000000000011110000100001000010101010110100111101011000101010110010100011;
        LUT[14] = 96'b110000001001000000000000000000000011110001001110110010000001100100111101100010110001000011011111;
        LUT[15] = 96'b110000001000100000000000000000000011110010000100110000011010011000111101101010100100010001010001;
        LUT[16] = 96'b110000001000000000000000000000000011110010101010011101100111000000111101110011111111100100011011;
        LUT[17] = 96'b110000000111000000000000000000000011110011011010111000001101110000111101111111010101110011100001;
        LUT[18] = 96'b110000000110000000000000000000000011110100001100100001011100111100111110000110011110000100100101;
        LUT[19] = 96'b110000000101000000000000000000000011110100110100011011110100100100111110001110100100111011011000;
        LUT[20] = 96'b110000000100000000000000000000000011110101100111101011101100100100111110011000001011111001111000;
        LUT[21] = 96'b110000000011000000000000000000000011110110010100101111100100011100111110100001101111110111111000;
        LUT[22] = 96'b110000000010000000000000000000000011110110111110111111010111101000111110101000010110010101111000;
        LUT[23] = 96'b110000000001000000000000000000000011110111110101001111000111011100111110101111111110100011100110;
        LUT[24] = 96'b110000000000000000000000000000000011111000011101011100011101101100111110111000101011110010000110;
        LUT[25] = 96'b101111111110000000000000000000000011111001001010001010011011111100111111000001001110111010110110;
        LUT[26] = 96'b101111111100000000000000000000000011111010000001110010101001000000111111000110100111011011111011;
        LUT[27] = 96'b101111111010000000000000000000000011111010100110101001111100000000111111001100011000000100111001;
        LUT[28] = 96'b101111111000000000000000000000000011111011010101111111010101011100111111010010010010110000000100;
        LUT[29] = 96'b101111110100000000000000000000000011111100001001011000100101000100111111010111111111011011000000;
        LUT[30] = 96'b101111110000000000000000000000000011111100110000011001111001010000111111011100110111100101100010;
        LUT[31] = 96'b101111101000000000000000000000000011111101100010100000100000110000111111100000000000000000000000;

        index = 0;
        
        valid_x_l = 1;
        
        reset = 1; 
        
        delay = 0;
        
        start_delaying = 0;
     end
 
    always @(posedge clock) begin
        if(compared) begin
            if(~x_lesser_than_x_l[0] && valid_x_l) begin
                if(reset) begin
                    valid_x_l = 0;
                    index = index + 10'b0000000001;
                    valid_x_l = 1;
                end
            end
            else begin
                valid_x_l = 0;
            end
            start_delaying = 1;    
        end
        if(start_delaying == 1) begin
            if(delay != 2'b10) begin
                reset = 0;
                delay = delay + 2'b01;
            end
            else begin
                reset = 1;
                delay = 0;
                start_delaying = 0;
            end
        end
    end
endmodule